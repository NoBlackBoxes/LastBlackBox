// AND Gate
module and_gate(Y, A, B);

  output Y;
  input A, B;

  assign Y = A & B;

endmodule
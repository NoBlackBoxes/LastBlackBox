// Hello World
module hello;

    // Initialize
    initial
        begin
            $display("Hello, World");
            $finish ;
        end

endmodule

// AND Gate
module and_gate(a, b, y);

    // Declarations
    input a;
    input b;
    output y;

    // Logic
    assign y = a & b;   // a AND b

endmodule
// ALU
module alu(src_A, src_B, ALU_control, ALU_result, zero);
    
    // Declarations
    input [31:0] src_A;
    input [31:0] src_B;
    input [2:0] ALU_control;
    output [31:0] ALU_result;
    output zero;

    // Intermediates

    // Logic

endmodule